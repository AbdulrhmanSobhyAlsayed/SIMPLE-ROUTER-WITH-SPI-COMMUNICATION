`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/26/2019 09:33:06 PM
// Design Name: 
// Module Name: SpiSlave
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
//
// Spi MODE 3: Output Edge: Falling, Data Capture: Rising
// MSB first data order
//
module SpiSlave(
    input sysClk,   // FPGA clock source
    input usrReset,
    //////////////////////////////////// 
    input  SCLK,    // Serial Clock: The clock pulses which synchronize data transmission generated by the master
    input  MOSI,    // SPI master out, slave in
    output MISO,   // SPI slave in, master out
    input  SS,     // SPI slave select
    ///////////////////////////////////
    output           rxValid,  // BYTE received is valid
	output reg [8:0] RX,       // BYTE received
	input [8:0]      TX);      // BYTE to transmit

    // Synchronize SCLK to FPGA clock using a two-stage shift-register
	// (bit [0] takes the hit of timing errors)
	reg [2:0] SCLKR;
	always @(posedge sysClk) 
	   SCLKR <= {SCLKR[1:0], SCLK};
	wire risingEdgeSCLK  = (SCLKR[2:1] == 2'b01);
	wire fallingEdgeSCLK = (SCLKR[2:1] == 2'b10);

    // Synchronize SS to FPGA clock using a two-stage shift-register
	reg [2:0] SSR;  
    always @(posedge sysClk) 
       SSR <= { SSR[1:0], SS };
	wire risingEdgeSS  = (SSR[2:1] == 2'b01);
	wire fallingEdgeSS = (SSR[2:1] == 2'b10);
	wire activeSS      = ~SSR[1];  // synchronous version of ~SS input
	       
	// Synchronize MOSI to FPGA clock using a two-stage shift-register
	reg [1:0] MOSIR;  
	always @(posedge sysClk) 
	   MOSIR <= { MOSIR[0], MOSI };
	wire syncMOSI = MOSIR[1];     // synchronous version of MOSI input    

    reg [3:0] byteCount;  // state corresponds to bit count
    reg MISOR = 1'bx;     //TX
    reg [8:0] data;      // Received data
    reg rxAvail = 1'b0;  // Reveived data is avaliable

    // next state logic
   wire [8:0] nextRX = {data[7:0], syncMOSI};
	
	// current state logic
	always @(posedge sysClk or posedge usrReset)
		if( usrReset )
			byteCount <= 4'd0;
		else  
		  if (activeSS)
            begin
			 if (fallingEdgeSS)  // begin of message
				byteCount <= 4'd0;
			 if (risingEdgeSCLK)  // bit available
				byteCount <= byteCount + 4'd1;
            end

	// output logic
	always @(posedge sysClk or posedge usrReset)
        if(usrReset)
        begin
            RX <= 9'hxx;
		    rxAvail <= 1'b0;
		end
		else
		  if (activeSS)  // Slave Select
            begin
                if (fallingEdgeSS)  // begin of message
                    rxAvail <= 1'b0;
                 // Receive
				if (risingEdgeSCLK)  // input on rising PCI clock edge (Data Capture [Received] on rising edge)
					if (byteCount == 4'd8) 
				    begin
					   RX <= nextRX;
					   rxAvail <= 1'b1;
				    end
					else
					begin
					   data <= nextRX;
					   rxAvail <= 1'b0;
					end
                   //Send
	            if (fallingEdgeSCLK)  // output on falling PCI clock edge (Data output [sent] on falling edge)
				    if (byteCount == 4'b000)
					begin 
					   data <= TX;  // load data with transmitted byte.
					   MISOR <= TX[8]; // Send the MSB 
				    end
				   else
					   MISOR <= data[8]; // Send the MSB
            end			
    
    assign MISO = activeSS ? MISOR : 1'bz;  // send MSB first
   // make rxAvail change on the falling edge, and make it 1 cycle wide
	reg rxAvailFall;
	reg rxAvailFallDelay;
	always @(negedge sysClk) 
	   rxAvailFall <= rxAvail;
	always @(negedge sysClk) 
	   rxAvailFallDelay <= rxAvailFall;
	assign rxValid = rxAvailFall & ~rxAvailFallDelay;            
endmodule
